`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date:    13:58:08 04/08/2017 
// Design Name: 
// Module Name:    testingsyntax 
// Project Name: 
// Target Devices: 
// Tool versions: 
// Description: 
//
// Dependencies: 
//
// Revision: 
// Revision 0.01 - File Created
// Additional Comments: 
//
//////////////////////////////////////////////////////////////////////////////////
module testingsyntax(a,b,c
    );
input [7:0]a;
input [7:0]b;
output [7:0]c;
assign c=a*b;


endmodule
